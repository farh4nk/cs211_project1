module toUpper_tb;

reg A0, A1, A2, A3, A4, A5, A6, A7;
wire B0, B1, B2, B3, B4, B5, B6, B7;

toUpper dut (.A0(A0), .A1(A1), .A2(A2), .A3(A3), .A4(A4), .A5(A5), .A6(A6), .A7(A7),
             .B0(B0), .B1(B1), .B2(B2), .B3(B3), .B4(B4), .B5(B5), .B6(B6), .B7(B7));

initial begin
    $dumpfile("toUpper.vcd");
    $dumpvars(0, toUpper_tb);
    
    // (
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00101000; #25;
    // H
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01001000; #25;
    // .
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10110111; #25;
    // f
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10000011; #25;
    // |
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111100; #25;
    // DC4
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00010100; #25;
    // ë
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b11101011; #25;
    // a
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01100001; #25;
    // A
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01000001; #25;
    // z
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111010; #25;
    // G
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01000111; #25;
    // m
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01101101; #25;
    // '
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10010010; #25;
    // 0
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00110000; #25;
    // Ï
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b11001111; #25;
    // : 
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00111010; #25;
    // {
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111011; #25;
    // ”
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10010100; #25;
    // DEL
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111111; #25;

    #50 $finish;
end

endmodule