`timescale 1ns / 1ps

module toUpper_tb;

reg A0, A1, A2, A3, A4, A5, A6, A7;
wire B0, B1, B2, B3, B4, B5, B6, B7;

toUpper dut (.A0(A0), .A1(A1), .A2(A2), .A3(A3), .A4(A4), .A5(A5), .A6(A6), .A7(A7),
             .B0(B0), .B1(B1), .B2(B2), .B3(B3), .B4(B4), .B5(B5), .B6(B6), .B7(B7));

initial begin
    $dumpfile("toUpper.vcd");
    $dumpvars(0, toUpper_tb);
    
    // (
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00101000; #10;
    // H
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01001000; #10;
    // .
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10110111; #10;
    // f
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10000011; #10;
    // |
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111100; #10;
    // DC4
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00010100; #10;
    // ë
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b11101011; #10;
    // a
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01100001; #10;
    // A
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01000001; #10;
    // z
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111010; #10;
    // G
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01000111; #10;
    // m
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01101101; #10;
    // '
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10010010; #10;
    // 0
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00110000; #10;
    // Ï
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b11001111; #10;
    // : 
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00111010; #10;
    // {
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111011; #10;
    // ”
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10010100; #10;
    // DEL
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111111; #10;

    #50 $finish;
end

endmodule