
module toUpper_tb;

reg A0, A1, A2, A3, A4, A5, A6, A7;
wire B0, B1, B2, B3, B4, B5, B6, B7;

toUpper dut (.A0(A0), .A1(A1), .A2(A2), .A3(A3), .A4(A4), .A5(A5), .A6(A6), .A7(A7),
             .B0(B0), .B1(B1), .B2(B2), .B3(B3), .B4(B4), .B5(B5), .B6(B6), .B7(B7));

initial begin
    $dumpfile("toUpper.vcd");
    $dumpvars(0, toUpper_tb);
    
    // (
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00101000; #15;
    // H
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01001000; #15;
    // .
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10110111; #15;
    // f
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10000011; #15;
    // |
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111100; #15;
    // DC4
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00010100; #15;
    // ë
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b11101011; #15;
    // a
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01100001; #15;
    // A
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01000001; #15;
    // z
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111010; #15;
    // G
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01000111; #15;
    // m
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01101101; #15;
    // '
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10010010; #15;
    // 0
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00110000; #15;
    // Ï
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b11001111; #15;
    // : 
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b00111010; #15;
    // {
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111011; #15;
    // ”
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b10010100; #15;
    // DEL
    {A7,A6,A5,A4,A3,A2,A1,A0} = 8'b01111111; #15;

    #50 $finish;
end

endmodule